module fix_decoder
#(

)
(

);

endmodule